module hex(input logic [15:0] in, output logic [7:0] out);

endmodule