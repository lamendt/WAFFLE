module UART(input logic clock,
input logic bitIn,
input logic [7:0] byteIn,
output logic bitOut,
output logic [7:0] byteOut);

endmodule
